/ictc/student_data/vantruong/final_pj/fn_prj_here/input_data/lef/RM_IHPSG13_1P_1024x16_c2_bm_bist.lef