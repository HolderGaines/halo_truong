/ictc/student_data/share/pd/data/user_setting/bondpad_70x70.lef