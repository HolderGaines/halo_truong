/ictc/student_data/vantruong/final_pj/fn_prj_here/input_data/lef/RM_IHPSG13_1P_4096x16_c3_bm_bist.lef