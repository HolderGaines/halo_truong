/ictc/student_data/vantruong/final_pj/fn_prj_here/input_data/lef/bondpad_70x70.lef