/ictc/student_data/vantruong/final_pj/fn_prj_here/input_data/lef/sg13g2_stdcell_weltap.lef