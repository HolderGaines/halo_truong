/ictc/student_data/share/pd/data/user_setting/sg13g2_io.lef